module rk_top(//
               rk_top_clk,rk_top_rst,rk_top_begin,MK_in,last,handshake,
               //
               rk,rk_top_addr,rk_top_en,rk_top_complete);

input rk_top_clk,rk_top_rst,rk_top_begin,last,handshake;
input[0:127] MK_in;


output rk_top_complete,rk_top_en;
output[0:4] rk_top_addr;
output[0:31] rk;

reg rk_top_complete,rk_top_en;
reg[0:4] rk_top_addr;
reg[0:5] currentstate,nextstate;    
reg[0:31] keyin1,keyin2,keyin3,keyin4,ck,rk;

wire[0:31] rkvar;
wire last,handshake;

reg aflag;
parameter  idle=6'b000000,
           ready=6'b000001,
           init=6'b000010,
           getrk1=6'b000011,
           getrk2=6'b000100,
           getrk3=6'b000101,
           getrk4=6'b000110,
           getrk5=6'b000111,
           getrk6=6'b001000,
           getrk7=6'b001001,
           getrk8=6'b001010,
           getrk9=6'b001011,
           getrk10=6'b001100,
           getrk11=6'b001101,
           getrk12=6'b001110,
           getrk13=6'b001111,
           getrk14=6'b010000,
           getrk15=6'b010001,
           getrk16=6'b010010,
           getrk17=6'b010011,
           getrk18=6'b010100,
           getrk19=6'b010101,
           getrk20=6'b010110,
           getrk21=6'b010111,
           getrk22=6'b011000,
           getrk23=6'b011001,
           getrk24=6'b011010,
           getrk25=6'b011011,
           getrk26=6'b011100,
           getrk27=6'b011101,
           getrk28=6'b011110,
           getrk29=6'b011111,
           getrk30=6'b100000,
           getrk31=6'b100001,
           getrk32=6'b100010,
           complete=6'b100011;

parameter FK0=32'h A3B1BAC6,FK1=32'h 56AA3350,FK2=32'h 677D9197,FK3=32'h b27022dc;

parameter CK0=32'h 00070e15, CK1=32'h 1c232a31, CK2=32'h 383f464d, CK3=32'h 545b6269,
          CK4=32'h 70777e85, CK5=32'h 8c939aa1, CK6=32'h a8afb6bd, CK7=32'h c4cbd2d9,
          CK8=32'h e0e7eef5, CK9=32'h fc030a11, CK10=32'h 181f262d,CK11=32'h 343b4249,
          CK12=32'h 50575e65,CK13=32'h 6c737a81,CK14=32'h 888f969d,CK15=32'h a4abb2b9,
          CK16=32'h c0c7ced5,CK17=32'h dce3eaf1,CK18=32'h f8ff060d,CK19=32'h 141b2229,
          CK20=32'h 30373e45,CK21=32'h 4c535a61,CK22=32'h 686f767d,CK23=32'h 848b9299,
          CK24=32'h a0a7aeb5,CK25=32'h bcc3cad1,CK26=32'h d8dfe6ed,CK27=32'h f4fb0209,
          CK28=32'h 10171e25,CK29=32'h 2c333a41,CK30=32'h 484f565d,CK31=32'h 646b7279;


always @(posedge rk_top_clk)
        if(~rk_top_rst||last)  
          begin		  
				currentstate<=idle;
			 end
        else
          currentstate<=nextstate; 



always @(currentstate or rk_top_begin or handshake)
        case(currentstate)
          idle:          begin                       
               if((rk_top_begin==1'b1)&&handshake)
                  begin
                 
                  	nextstate<=ready;
		  end
               else
                  nextstate<=idle;  					
						end
          ready:                                
               if((rk_top_begin==1'b1)&&handshake)
                  begin
                  	nextstate<=init;
		  end
               else
                  nextstate<=idle;
          init:                                
               nextstate<=getrk1;
          getrk1:
               nextstate<=getrk2;             
          getrk2:
               nextstate<=getrk3;
          getrk3:
               nextstate<=getrk4;
          getrk4:
               nextstate<=getrk5;
          getrk5:
               nextstate<=getrk6;
          getrk6:
               nextstate<=getrk7;
          getrk7:
               nextstate<=getrk8;
          getrk8:
               nextstate<=getrk9;
          getrk9:
               nextstate<=getrk10;
          getrk10:
               nextstate<=getrk11;
          getrk11:
               nextstate<=getrk12;     
          getrk12:
               nextstate<=getrk13;
          getrk13:
               nextstate<=getrk14;
          getrk14:
               nextstate<=getrk15;
          getrk15:
               nextstate<=getrk16;
          getrk16:
               nextstate<=getrk17;
          getrk17:
               nextstate<=getrk18;
          getrk18:
               nextstate<=getrk19;
          getrk19:
               nextstate<=getrk20;
          getrk20:
               nextstate<=getrk21;
          getrk21:
               nextstate<=getrk22;     
          getrk22:
               nextstate<=getrk23;
          getrk23:
               nextstate<=getrk24;
          getrk24:
               nextstate<=getrk25;
          getrk25:
               nextstate<=getrk26;
          getrk26:
               nextstate<=getrk27;
          getrk27:
               nextstate<=getrk28;
          getrk28:
               nextstate<=getrk29;
          getrk29:
               nextstate<=getrk30;
          getrk30:
               nextstate<=getrk31;
          getrk31:
               nextstate<=getrk32;
          getrk32:
               nextstate<=complete;
          complete:
               nextstate<=idle;
          default:
               nextstate<=idle;
        endcase

//״̬ʵֵĹܡ
always @(posedge rk_top_clk)
        case(nextstate)
          idle:                                             
               begin
                  rk<=32'bz; 
						if(last) 
						rk_top_complete<=1'b0;
						
               end
          ready:                                           
               begin
 		            rk_top_en<=1'b0;
                  rk_top_addr<=5'b00000;
                  rk<=32'bz;
                  keyin1<=MK_in[0:31];
                  keyin2<=MK_in[32:63];
                  keyin3<=MK_in[64:95];   
                  keyin4<=MK_in[96:127];
               end
          init:                                            
               begin
                  ck<=CK0;
						rk_top_complete<=1'b0;
                  keyin1<=keyin1^FK0;
                  keyin2<=keyin2^FK1;
                  keyin3<=keyin3^FK2;   
                  keyin4<=keyin4^FK3;
               end
          getrk1:                                          
               begin
                  rk_top_en<=1'b1;
                  rk<=rkvar;
                  ck<=CK1;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk2:                                         
               begin
                  rk_top_addr<=5'b00001;
                  rk<=rkvar;
                  ck<=CK2;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk3:
               begin
                  rk_top_addr<=5'b00010;
                  rk<=rkvar;
                  ck<=CK3;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk4:
               begin
                  rk_top_addr<=5'b00011;
                  rk<=rkvar;
                  ck<=CK4;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk5:
               begin
                  rk_top_addr<=5'b00100;
                  rk<=rkvar;
                  ck<=CK5;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk6:
               begin
                  rk_top_addr<=5'b00101;
                  rk<=rkvar;
                  ck<=CK6;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk7:
               begin
                  rk_top_addr<=5'b00110;
                  rk<=rkvar;
                  ck<=CK7;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk8:
               begin
                  rk_top_addr<=5'b00111;
                  rk<=rkvar;
                  ck<=CK8;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk9:
               begin
                  rk_top_addr<=5'b01000;
                  rk<=rkvar;
                  ck<=CK9;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk10:
               begin
                  rk_top_addr<=5'b01001;
                  rk<=rkvar;
                  ck<=CK10;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk11:
               begin
                  rk_top_addr<=5'b01010;
                  rk<=rkvar;
                  ck<=CK11;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end     
          getrk12:
               begin
                  rk_top_addr<=5'b01011;
                  rk<=rkvar;
                  ck<=CK12;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk13:
               begin
                  rk_top_addr<=5'b01100;
                  rk<=rkvar;
                  ck<=CK13;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk14:
               begin
                  rk_top_addr<=5'b01101;
                  rk<=rkvar;
                  ck<=CK14;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk15:
               begin
                  rk_top_addr<=5'b01110;
                  rk<=rkvar;
                  ck<=CK15;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk16:
               begin
                  rk_top_addr<=5'b01111;
                  rk<=rkvar;
                  ck<=CK16;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk17:
               begin
                  rk_top_addr<=5'b10000;
                  rk<=rkvar;
                  ck<=CK17;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk18:
               begin
                  rk_top_addr<=5'b10001;
                  rk<=rkvar;
                  ck<=CK18;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk19:
               begin
                  rk_top_addr<=5'b10010;
                  rk<=rkvar;
                  ck<=CK19;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk20:
               begin
                  rk_top_addr<=5'b10011;
                  rk<=rkvar;
                  ck<=CK20;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk21:
               begin
                  rk_top_addr<=5'b10100;
                  rk<=rkvar;
                  ck<=CK21;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end     
          getrk22:
               begin
                  rk_top_addr<=5'b10101;
                  rk<=rkvar;
                  ck<=CK22;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk23:
               begin
                  rk_top_addr<=5'b10110;
                  rk<=rkvar;
                  ck<=CK23;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk24:
               begin
                  rk_top_addr<=5'b10111;
                  rk<=rkvar;
                  ck<=CK24;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk25:
               begin
                  rk_top_addr<=5'b11000;
                  rk<=rkvar;
                  ck<=CK25;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk26:
               begin
                  rk_top_addr<=5'b11001;
                  rk<=rkvar;
                  ck<=CK26;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk27:
               begin
                  rk_top_addr<=5'b11010;
                  rk<=rkvar;
                  ck<=CK27;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk28:
               begin
                  rk_top_addr<=5'b11011;
                  rk<=rkvar;
                  ck<=CK28;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk29:
               begin
                  rk_top_addr<=5'b11100;
                  rk<=rkvar;
                  ck<=CK29;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk30:
               begin
                  rk_top_addr<=5'b11101;
                  rk<=rkvar;
                  ck<=CK30;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk31:
               begin
                  rk_top_addr<=5'b11110;
                  rk<=rkvar;
                  ck<=CK31;
                  keyin1<=keyin2;
                  keyin2<=keyin3;
                  keyin3<=keyin4;
                  keyin4<=rkvar;
               end
          getrk32:
               begin
                  rk_top_addr<=5'b11111;
                  rk<=rkvar;
               end
          complete:
               begin
                  rk_top_en<=1'b0;
                  rk_top_complete<=1'b1;               
               end
          default:
               begin
                  rk_top_complete<=1'b0;
                  rk_top_en<=1'b0;
                  rk_top_addr<=5'b00000;
                  rk<=32'bz; 
               end
      endcase            

Frk_function Frk_rk_top(keyin1,keyin2,keyin3,keyin4,ck,rkvar);  
    
endmodule	